`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:47:36 12/03/2017 
// Design Name: 
// Module Name:    ctrl 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ctrl(
    input  [31:0] Instr,
    input  Branch,
	 input  INT_REQ,
    output Mem_Write,
    output Reg_Write,
    output [3:0] ALU_Op,
    output Shift,
	 output EXT_Op,
    output ALU_B_Sel,
    output [2:0] PC_Src,
    output [1:0] Data_To_Reg,
    output [1:0] Reg_Dst,
	 output OP_EXP,
	 output [1:0] WT_PR
    );
	 wire [5:0] Op		= Instr[31:26];
	 wire [5:0] Func	= Instr[5:0];
	 wire [4:0] Id		= Instr[20:16];
	 wire [4:0] Wt		= Instr[25:21];
	 wire [18:0] control;
	 
	 assign {WT_PR,OP_EXP,Mem_Write,Reg_Write,ALU_Op,Shift,ALU_B_Sel, EXT_Op, PC_Src, Data_To_Reg, Reg_Dst} = control;
	 assign control =
			(INT_REQ)			? 19'b00_0_0_0_0000_0_0_0_100_00_00 : //Interrupt
			(Op == 6'b100011) ? 19'b00_0_0_1_0000_0_1_1_000_01_00 : //lw
			(Op == 6'b100000) ? 19'b00_0_0_1_0000_0_1_1_000_01_00 : //lb
			(Op == 6'b100100) ? 19'b00_0_0_1_0000_0_1_1_000_01_00 : //lbu
			(Op == 6'b100001) ? 19'b00_0_0_1_0000_0_1_1_000_01_00 : //lh
			(Op == 6'b100101) ? 19'b00_0_0_1_0000_0_1_1_000_01_00 : //lhu
			(Op == 6'b101011) ? 19'b00_0_1_0_0000_0_1_1_000_00_00 : //sw
			(Op == 6'b101000) ? 19'b00_0_1_0_0000_0_1_1_000_00_00 : //sb
			(Op == 6'b101001) ? 19'b00_0_1_0_0000_0_1_1_000_00_00 : //sh
			
			
			(Op == 6'b000100 || Op == 6'b000101 || Op == 6'b000111 || Op == 6'b000110) ? ((Branch) ? 19'b00_0_0_0_0100_0_0_1_001_00_00 : 19'b00_0_0_0_0100_0_0_1_000_00_00) : //beq bne bgtz blez

			(Op == 6'b000001 && (Id == 5'b00000 || Id == 5'b00001)) ? ((Branch) ? 19'b00_0_0_0_0100_0_0_1_001_00_00 : 19'b00_0_0_0_0100_0_0_1_000_00_00) : //bgez bltz
			
			(Op == 6'b000001 && !(Id == 5'b00000 || Id == 5'b00001)) ? ((Branch) ? 19'b00_0_0_1_0100_0_0_1_001_10_10 : 19'b00_0_0_0_0100_0_0_1_000_10_10) : //bgezal bltzal
	
					
			(Op == 6'b000010) ? 19'b00_0_0_0_0000_0_0_0_011_00_00 : //j
			(Op == 6'b000011) ? 19'b00_0_0_1_0000_0_0_0_011_10_10 : //jal
			
			
			(Op == 6'b001111) ? 19'b00_0_0_1_0110_0_1_0_000_00_00 : //lui
			(Op == 6'b001000) ? 19'b00_0_0_1_1001_0_1_1_000_00_00 : //addi
			(Op == 6'b001001) ? 19'b00_0_0_1_0000_0_1_1_000_00_00 : //addiu
			(Op == 6'b001100) ? 19'b00_0_0_1_0001_0_1_0_000_00_00 : //andi
			(Op == 6'b001101) ? 19'b00_0_0_1_0101_0_1_0_000_00_00 : //ori
			(Op == 6'b001110) ? 19'b00_0_0_1_0010_0_1_0_000_00_00 : //xori
			
			(Op == 6'b001010) ? 19'b00_0_0_1_0100_0_1_1_000_00_00 : //slti
		   (Op == 6'b001011) ? 19'b00_0_0_1_1000_0_1_1_000_00_00 : //sltiu

			//COP0
			(Op == 6'b010000 && Wt == 5'b00000) ? 19'b10_0_0_1_0000_0_0_0_000_01_00 : //mfc0
			(Op == 6'b010000 && Wt == 5'b00100) ? 19'b01_0_0_0_0000_0_0_0_000_00_01 : //mtc0
			(Op == 6'b010000 && Wt == 5'b10000) ? 19'b11_0_0_0_0000_0_0_0_101_00_00 : //eret
				 
			(Op == 6'b000000) ? //R
					  ((Func == 6'b100000) ? 19'b00_0_0_1_1001_0_0_0_000_00_01 : //add
						(Func == 6'b100001) ? 19'b00_0_0_1_0000_0_0_0_000_00_01 : //addu
						(Func == 6'b100010) ? 19'b00_0_0_1_0100_0_0_0_000_00_01 : //sub
						(Func == 6'b100011) ? 19'b00_0_0_1_1000_0_0_0_000_00_01 : //subu
						(Func == 6'b100100) ? 19'b00_0_0_1_0001_0_0_0_000_00_01 : //and
						(Func == 6'b100101) ? 19'b00_0_0_1_0101_0_0_0_000_00_01 : //or
						(Func == 6'b100110) ? 19'b00_0_0_1_0010_0_0_0_000_00_01 : //xor						
						(Func == 6'b100111) ? 19'b00_0_0_1_1110_0_0_0_000_00_01 : //nor
						
						
						(Func == 6'b000010) ? 19'b00_0_0_1_0111_1_0_0_000_00_01 : //srl
						(Func == 6'b000011) ? 19'b00_0_0_1_1111_1_0_0_000_00_01 : //sra
						(Func == 6'b000100) ? 19'b00_0_0_1_0011_0_0_0_000_00_01 : //sllv
						(Func == 6'b000110) ? 19'b00_0_0_1_0111_0_0_0_000_00_01 : //srlv
						(Func == 6'b000111) ? 19'b00_0_0_1_1111_0_0_0_000_00_01 : //srav
						
						(Func == 6'b001000) ? 19'b00_0_0_0_0000_0_0_0_010_00_00 : //jr
						(Func == 6'b001001) ? 19'b00_0_0_1_0000_0_0_0_010_10_01 : //jalr
						
						
						(Func == 6'b101010) ? 19'b00_0_0_1_0100_0_0_0_000_00_01 : //slt
						(Func == 6'b101011) ? 19'b00_0_0_1_1000_0_0_0_000_00_01 : //sltu
						
						
						(Func == 6'b011010) ? 19'b00_0_0_0_0000_0_0_0_000_00_00 : //div
						(Func == 6'b011011) ? 19'b00_0_0_0_0000_0_0_0_000_00_00 : //divu
						(Func == 6'b011000) ? 19'b00_0_0_0_0000_0_0_0_000_00_00 : //mult
						(Func == 6'b011001) ? 19'b00_0_0_0_0000_0_0_0_000_00_00 : //multu
						(Func == 6'b010000) ? 19'b00_0_0_1_0000_0_0_0_000_00_01 : //mfhi
						(Func == 6'b010010) ? 19'b00_0_0_1_0000_0_0_0_000_00_01 : //mflo
						(Func == 6'b010001) ? 19'b00_0_0_0_0000_0_0_0_000_00_00 : //mthi
						(Func == 6'b010011) ? 19'b00_0_0_0_0000_0_0_0_000_00_00 : //mtlo
						(Func == 6'b000000) ? ((Instr == 32'b0) ? 19'b00_0_0_0_0000_0_0_0_000_00_00 : 19'b00_0_0_1_0011_1_0_0_000_00_01) : 19'b01_1_0_0_0000_0_0_0_000_00_00) : //nop sll
													 19'b01_1_0_0_0000_0_0_0_000_00_00 ;
endmodule
